library IEEE;
use IEEE.std_logic_1164.all;

entity Mux_tb is
end;

architecture Mux_tb_arq of Mux_tb is
    -- Parte declarativa
    component Mux is
        port(
            a_i: in std_logic;
			b_i: in std_logic;
			sel_i: in std_logic;
			s_o: out std_logic
        );
    end component;

    -- Declaracion de senales de prueba
	signal a_tb: std_logic := '0';
	signal b_tb: std_logic := '1';
	signal sel_tb: std_logic := '0';
	signal s_tb: std_logic;

begin 

    -- a_tb <= '1' after 100 ns, '0' after 500 ns;
	-- b_tb <= '1' after 200 ns, '0' after 400 ns;
	-- ci_tb <= '1' after 150 ns, '0' after 900 ns;
	a_tb <= '1' after 100 ns;
	b_tb <= '0' after 70 ns;
	sel_tb <= '1' after 40 ns, '0' after 130 ns;

    DUT: Mux
    port map(
            a_i	 => a_tb, 
			b_i	 => b_tb,
			sel_i => sel_tb,
			s_o	 => s_tb
    );
end;