library IEEE;
use IEEE.std_logic_1164.all;

entity comp is
    port(
        a_i : in std_logic;
        s_o : out std_logic
    );
end;

architecture comp_arq of comp is
    -- Parte declarativa
begin   
    -- Parte descriptiva
end;